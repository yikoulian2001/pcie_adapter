
parameter	DWIDTH = 256;
parameter	MAXTAG = 64;

static bit[7:0] MEMORY[bit[63:0]];
